//created by jiemin on 20150909
//asynchronous fifo -- systemverilog testbench
module tb;

endmodule
