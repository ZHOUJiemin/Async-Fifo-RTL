//created by jiemin on 20150910
//asynchronous fifo -- test program class Scoreboard
class Scoreboard;

endclass
